module SPI_driver (
    input logic clk,
    input logic rst,
    input logic [7:0] data_in,
    input logic SPI_MISO, // Slave Out (Master In)
    input logic SPI_start,
    output logic SPI_MOSI, // Master Out (Slave In)
    output logic SPI_CLK,
    output logic SPI_EN, // Slave Select (SS)
    output logic [7:0] data_out
);

// State definitions
typedef enum {
    IDLE,
    SEND,
    RECEIVE
} state_t;

state_t state = IDLE;

// Internal signals
logic [7:0] tx_data;
logic [7:0] rx_data;
logic [2:0] bit_count;
logic [1:0] cpol_ch;

// Edge detection for clock
logic clk_prev = 0;

// CPOL and CPHA settings
// CPOL=1 (Idle high), CPHA=1 (Sample on rising edge)
assign cpol_ch = 2'b11;

// Initializing variables
initial begin
    tx_data = 0;
    rx_data = 0;
end

always_ff @(posedge clk) begin
    if (rst) begin
        state <= IDLE;
        tx_data <= 0;
        rx_data <= 0;
        bit_count <= 0;
        SPI_MOSI <= 0;
        SPI_CLK <= 1; // Idle high
        SPI_EN <= 1;  // SS high (not selected)
        data_out <= 0;
        clk_prev <= 0;
    end else begin
        // Clock generation logic
        if (state == SEND || state == RECEIVE) begin
            // Generate clock based on CPOL and CPHA
            if (bit_count < 8) begin
                // Toggle clock
                SPI_CLK <= ~SPI_CLK;
            end
        end
        
        // Edge detection
        if (clk != clk_prev) begin
            // Rising edge detection
            if (SPI_CLK && !clk_prev) begin
                // Data capture on rising edge for receiving
                if (state == RECEIVE) begin
                    rx_data <= {rx_data[6:0], SPI_MISO};
                end
            end
        end
        
        case (state)
            IDLE: begin
                if (SPI_start) begin
                    // Select slave (SS) by driving low
                    SPI_EN <= 0;
                    state <= SEND;
                    tx_data <= data_in;
                    bit_count <= 0;
                    // Send first bit (MSB)
                    SPI_MOSI <= (tx_data >> (7 - bit_count)) & 1;
                    bit_count <= bit_count + 1;
                end
            end
            
            SEND: begin
                if (bit_count < 8) begin
                    // Shift out data on rising edge
                    SPI_MOSI <= (tx_data >> (7 - bit_count)) & 1;
                    // Toggle clock
                    bit_count <= bit_count + 1;
                    
                    if (bit_count == 8) begin
                        // Last bit sent
                        SPI_CLK <= 1; // Ensure clock stops
                        // If there's data to receive, switch to receive state
                        if (data_in == 0) begin
                            state <= RECEIVE;
                            rx_data <= 0;
                            bit_count <= 0;
                        end else begin
                            // No data to receive, return to idle
                            state <= IDLE;
                            SPI_EN <= 1; // Deselect
                        end
                    end
                end
            end
            
            RECEIVE: begin
                if (bit_count < 8) begin
                    // On the rising edge, data is captured
                    rx_data <= {rx_data[6:0], SPI_MISO};
                    bit_count <= bit_count + 1;
                    
                    if (bit_count == 8) begin
                        data_out <= rx_data;
                        state <= IDLE;
                        // Deselect slave
                        SPI_EN <= 1;
                    end
                end
            end
        endcase
        
        clk_prev <= clk;
    end
end

// Immediate output assignments for non-stateful signals (should be moved into the always_ff block above)
assign SPI_CLK = 1; // To be generated by the state machine

endmodule