// -----------------------------------------------------------------------------
// Simple 8-bit SPI Master (Mode-2 : CPOL = 1, CPHA = 0)
// ‑ CPOL = 1 : SCLK is HIGH when bus is idle
// ‑ CPHA = 0 : Data is driven valid before the first (falling) edge;
//              data is captured on the first (falling) edge.
//
// Generic, single-byte transaction started with SPI_start.
// Clock is generated by dividing the system clock (clk) by parameter CLK_DIV*2.
// -----------------------------------------------------------------------------
module SPI_driver #(
    parameter int unsigned CLK_DIV = 4   // sys_clk ticks per half SCLK period
)(
    input  logic        clk,        // system clock
    input  logic        rst,        // synchronous, active high reset
    input  logic [7:0]  data_in,    // byte to be transmitted
    input  logic        SPI_MISO,   // slave -> master data
    input  logic        SPI_start,  // assert for one clk to start transfer
    output logic        SPI_MOSI,   // master -> slave data
    output logic        SPI_CLK,    // serial clock (CPOL = 1)
    output logic        SPI_EN,     // chip-select (active low)
    output logic [7:0]  data_out    // byte just received
);

    // ---------------------------------------------------------
    // Local registers / signals
    // ---------------------------------------------------------
    typedef enum logic [1:0] {IDLE, ASSERT_CS, TRANSFER, DEASSERT_CS} state_t;
    state_t          state, nxt_state;

    logic [$clog2(CLK_DIV)-1:0] clk_cnt;   // clock divider counter
    logic                        sclk_int; // internal clock (pre-CPOL ORed)
    logic [7:0]                  shreg;    // shift register (Tx/Rx)
    logic [2:0]                  bit_cnt;  // tracks 0->7
    logic                        sclk_fall;// single-cycle pulse – SCLK falling
    logic                        sclk_rise;// single-cycle pulse – SCLK rising

    // ---------------------------------------------------------
    // Clock divider – produces sclk_int toggles
    // ---------------------------------------------------------
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            clk_cnt  <= '0;
            sclk_int <= 1'b0;
        end
        else if (state == TRANSFER) begin
            if (clk_cnt == CLK_DIV-1) begin
                clk_cnt  <= '0;
                sclk_int <= ~sclk_int;
            end
            else begin
                clk_cnt <= clk_cnt + 1'b1;
            end
        end
        else begin
            clk_cnt  <= '0;
            sclk_int <= 1'b0;   // ensure defined after IDLE
        end
    end

    // Create single-cycle edge indicators
    logic sclk_int_d;
    always_ff @(posedge clk) sclk_int_d <= sclk_int;
    assign sclk_rise =  sclk_int & ~sclk_int_d;
    assign sclk_fall = ~sclk_int &  sclk_int_d;

    // ---------------------------------------------------------
    // Main FSM
    // ---------------------------------------------------------
    always_ff @(posedge clk or posedge rst) begin
        if (rst) state <= IDLE;
        else     state <= nxt_state;
    end

    always_comb begin
        nxt_state = state;
        case (state)
            IDLE        : if (SPI_start)      nxt_state = ASSERT_CS;
            ASSERT_CS   :                    nxt_state = TRANSFER;
            TRANSFER    : if (bit_cnt == 3'd7 && sclk_rise)
                                               nxt_state = DEASSERT_CS;
            DEASSERT_CS :                    nxt_state = IDLE;
        endcase
    end

    // ---------------------------------------------------------
    // Bit counter
    // ---------------------------------------------------------
    always_ff @(posedge clk or posedge rst) begin
        if (rst) bit_cnt <= 3'd0;
        else if (state == ASSERT_CS)  bit_cnt <= 3'd0;
        else if (state == TRANSFER && sclk_rise)
            bit_cnt <= bit_cnt + 1'b1;
    end

    // ---------------------------------------------------------
    // Shift register – CPOL=1, CPHA=0 protocol handling
    //  • MOSI must be valid before the falling edge.
    //  • MISO is sampled on the falling edge.
    // ---------------------------------------------------------
    // Load on ASSERT_CS
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            shreg <= 8'h00;
        end
        else begin
            case (state)
                ASSERT_CS : shreg <= data_in;         // load Tx data
                TRANSFER  : begin
                    // Falling edge : sample MISO into LSB
                    if (sclk_fall)
                        shreg <= {shreg[6:0], SPI_MISO};
                    // Rising edge  : shift for next bit
                    if (sclk_rise)
                        shreg <= {shreg[6:0], 1'b0};
                end
            endcase
        end
    end

    // ---------------------------------------------------------
    // Outputs
    // ---------------------------------------------------------
    // SCLK : CPOL=1 -> idle HIGH
    assign SPI_CLK = (state == TRANSFER) ? ~sclk_int : 1'b1; // invert to get falling first edge

    // MOSI is always the current MSB (bit 7) of shift register
    always_ff @(posedge clk or posedge rst) begin
        if (rst)            SPI_MOSI <= 1'b0;
        // update before next falling edge (i.e. after rising edge shift)
        else if (state == ASSERT_CS)        SPI_MOSI <= shreg[7];
        else if (state == TRANSFER && sclk_rise)
                                SPI_MOSI <= shreg[7];
    end

    // Chip-select (active low)
    assign SPI_EN = (state == TRANSFER || state == ASSERT_CS) ? 1'b0 : 1'b1;

    // Present captured byte once transfer is complete
    always_ff @(posedge clk or posedge rst) begin
        if (rst)                   data_out <= 8'h00;
        else if (state == DEASSERT_CS) data_out <= shreg;
    end

endmodule